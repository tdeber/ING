module EJ1(
    input wire A,
    input wire B,
    output wire X
);

// Operación lógica AND entre A y B
assign X = A & B;

endmodule

