`include "Sumador/suma.v"
module alu(
     input wire In1,In2,CBin,
     input wire [2:0] cod,
     output wire Rta,CBout
    );
    //Necesito hacer un case y para cada opcion llamo al modulo q le corresponde
    


endmodule
